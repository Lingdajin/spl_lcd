// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.13.0.56.2
// Netlist written on Wed Jan 15 19:58:40 2025
//
// Verilog Description of module rom_8x4096
//

module rom_8x4096 (Address, OutClock, OutClockEn, Reset, Q) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(8[8:18])
    input [11:0]Address;   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    input OutClock;   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(10[16:24])
    input OutClockEn;   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(11[16:26])
    input Reset;   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(12[16:21])
    output [7:0]Q;   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    
    wire OutClock_c /* synthesis is_clock=1 */ ;   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(10[16:24])
    
    wire Address_c_11, Address_c_10, Address_c_9, Address_c_8, Address_c_7, 
        Address_c_6, Address_c_5, Address_c_4, Address_c_3, Address_c_2, 
        Address_c_1, Address_c_0, OutClockEn_c, Reset_c, Q_c_7, Q_c_6, 
        Q_c_5, Q_c_4, Q_c_3, Q_c_2, Q_c_1, Q_c_0, scuba_vlo, VCC_net;
    
    OB Q_pad_2 (.I(Q_c_2), .O(Q[2]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    OB Q_pad_3 (.I(Q_c_3), .O(Q[3]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    OB Q_pad_4 (.I(Q_c_4), .O(Q[4]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    DP8KC rom_8x4096_0_3_0 (.DIA0(scuba_vlo), .DIA1(scuba_vlo), .DIA2(scuba_vlo), 
          .DIA3(scuba_vlo), .DIA4(scuba_vlo), .DIA5(scuba_vlo), .DIA6(scuba_vlo), 
          .DIA7(scuba_vlo), .DIA8(scuba_vlo), .ADA0(scuba_vlo), .ADA1(Address_c_0), 
          .ADA2(Address_c_1), .ADA3(Address_c_2), .ADA4(Address_c_3), 
          .ADA5(Address_c_4), .ADA6(Address_c_5), .ADA7(Address_c_6), 
          .ADA8(Address_c_7), .ADA9(Address_c_8), .ADA10(Address_c_9), 
          .ADA11(Address_c_10), .ADA12(Address_c_11), .CEA(OutClockEn_c), 
          .OCEA(OutClockEn_c), .CLKA(OutClock_c), .WEA(scuba_vlo), .CSA0(scuba_vlo), 
          .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(Reset_c), .DIB0(scuba_vlo), 
          .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
          .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
          .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), .ADB3(scuba_vlo), 
          .ADB4(scuba_vlo), .ADB5(scuba_vlo), .ADB6(scuba_vlo), .ADB7(scuba_vlo), 
          .ADB8(scuba_vlo), .ADB9(scuba_vlo), .ADB10(scuba_vlo), .ADB11(scuba_vlo), 
          .ADB12(scuba_vlo), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(scuba_vlo), 
          .WEB(scuba_vlo), .CSB0(scuba_vlo), .CSB1(scuba_vlo), .CSB2(scuba_vlo), 
          .RSTB(scuba_vlo), .DOA0(Q_c_6), .DOA1(Q_c_7)) /* synthesis MEM_LPC_FILE="rom_8x4096.lpc", MEM_INIT_FILE="rom_8x4096.mem", syn_instantiated=1 */ ;
    defparam rom_8x4096_0_3_0.DATA_WIDTH_A = 2;
    defparam rom_8x4096_0_3_0.DATA_WIDTH_B = 2;
    defparam rom_8x4096_0_3_0.REGMODE_A = "NOREG";
    defparam rom_8x4096_0_3_0.REGMODE_B = "NOREG";
    defparam rom_8x4096_0_3_0.CSDECODE_A = "0b000";
    defparam rom_8x4096_0_3_0.CSDECODE_B = "0b111";
    defparam rom_8x4096_0_3_0.WRITEMODE_A = "NORMAL";
    defparam rom_8x4096_0_3_0.WRITEMODE_B = "NORMAL";
    defparam rom_8x4096_0_3_0.GSR = "ENABLED";
    defparam rom_8x4096_0_3_0.RESETMODE = "ASYNC";
    defparam rom_8x4096_0_3_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam rom_8x4096_0_3_0.INIT_DATA = "STATIC";
    defparam rom_8x4096_0_3_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_09 = "0x0000000800000000000600200000010A800000000000000000020100000000000028000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_0A = "0x0AA5400000000010C000000000000000600000000000000000002000000000810000000000000010";
    defparam rom_8x4096_0_3_0.INITVAL_0B = "0x0A0150000000000080000A800000000A8000800402000000000A8050000500015000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_0C = "0x08A54000000005500000002000000002010000040000008000000000000000000000000AA5400001";
    defparam rom_8x4096_0_3_0.INITVAL_0D = "0x0AA55180000080000000000010000108001000000AA540000008005080000A8000000D0800000000";
    defparam rom_8x4096_0_3_0.INITVAL_0E = "0x00055000000AA54000050AA55180040000008005000000000400000080000000008000000000000D";
    defparam rom_8x4096_0_3_0.INITVAL_0F = "0x000011800000A550800000005180010AA551800000001080010A0050800D00015000100AA5400000";
    defparam rom_8x4096_0_3_0.INITVAL_10 = "0x00000000C0000000000000000020000000000050000000001000000008010800008000000000800D";
    defparam rom_8x4096_0_3_0.INITVAL_11 = "0x0AA00000140004000000000421800100A000000D0AA550800100200000000A8000000D0AA0000000";
    defparam rom_8x4096_0_3_0.INITVAL_12 = "0x0A800000010AA000000D0AA000000A1544000000000000000400040000000000000000000000000D";
    defparam rom_8x4096_0_3_0.INITVAL_13 = "0x00040000000AAC000000002C00000D0AA40000000000000001082400000000240000D50AA4000000";
    defparam rom_8x4096_0_3_0.INITVAL_14 = "0x0000000000000000000000000060000000000000000000003000000018050004000000002C000004";
    defparam rom_8x4096_0_3_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_3_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    OB Q_pad_5 (.I(Q_c_5), .O(Q[5]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    OB Q_pad_6 (.I(Q_c_6), .O(Q[6]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    DP8KC rom_8x4096_0_0_3 (.DIA0(scuba_vlo), .DIA1(scuba_vlo), .DIA2(scuba_vlo), 
          .DIA3(scuba_vlo), .DIA4(scuba_vlo), .DIA5(scuba_vlo), .DIA6(scuba_vlo), 
          .DIA7(scuba_vlo), .DIA8(scuba_vlo), .ADA0(scuba_vlo), .ADA1(Address_c_0), 
          .ADA2(Address_c_1), .ADA3(Address_c_2), .ADA4(Address_c_3), 
          .ADA5(Address_c_4), .ADA6(Address_c_5), .ADA7(Address_c_6), 
          .ADA8(Address_c_7), .ADA9(Address_c_8), .ADA10(Address_c_9), 
          .ADA11(Address_c_10), .ADA12(Address_c_11), .CEA(OutClockEn_c), 
          .OCEA(OutClockEn_c), .CLKA(OutClock_c), .WEA(scuba_vlo), .CSA0(scuba_vlo), 
          .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(Reset_c), .DIB0(scuba_vlo), 
          .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
          .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
          .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), .ADB3(scuba_vlo), 
          .ADB4(scuba_vlo), .ADB5(scuba_vlo), .ADB6(scuba_vlo), .ADB7(scuba_vlo), 
          .ADB8(scuba_vlo), .ADB9(scuba_vlo), .ADB10(scuba_vlo), .ADB11(scuba_vlo), 
          .ADB12(scuba_vlo), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(scuba_vlo), 
          .WEB(scuba_vlo), .CSB0(scuba_vlo), .CSB1(scuba_vlo), .CSB2(scuba_vlo), 
          .RSTB(scuba_vlo), .DOA0(Q_c_0), .DOA1(Q_c_1)) /* synthesis MEM_LPC_FILE="rom_8x4096.lpc", MEM_INIT_FILE="rom_8x4096.mem", syn_instantiated=1 */ ;
    defparam rom_8x4096_0_0_3.DATA_WIDTH_A = 2;
    defparam rom_8x4096_0_0_3.DATA_WIDTH_B = 2;
    defparam rom_8x4096_0_0_3.REGMODE_A = "NOREG";
    defparam rom_8x4096_0_0_3.REGMODE_B = "NOREG";
    defparam rom_8x4096_0_0_3.CSDECODE_A = "0b000";
    defparam rom_8x4096_0_0_3.CSDECODE_B = "0b111";
    defparam rom_8x4096_0_0_3.WRITEMODE_A = "NORMAL";
    defparam rom_8x4096_0_0_3.WRITEMODE_B = "NORMAL";
    defparam rom_8x4096_0_0_3.GSR = "ENABLED";
    defparam rom_8x4096_0_0_3.RESETMODE = "ASYNC";
    defparam rom_8x4096_0_0_3.ASYNC_RESET_RELEASE = "SYNC";
    defparam rom_8x4096_0_0_3.INIT_DATA = "STATIC";
    defparam rom_8x4096_0_0_3.INITVAL_00 = "0x0D200040000100000000000000D0090B480014090C00D01260014E300000000A0000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_01 = "0x0E00013400012000C00D1026001000100090AA600348000008000000000C00068000000000C00000";
    defparam rom_8x4096_0_0_3.INITVAL_02 = "0x000010C00800008000C30000001000000000000000000014250C0090B260000000E0090BA600120D";
    defparam rom_8x4096_0_0_3.INITVAL_03 = "0x00020018000600E154B0004551000E154B001CAA1600E154B0012550C00E154B001CA8000090AA60";
    defparam rom_8x4096_0_0_3.INITVAL_04 = "0x160080007001A090C00E154B0012D50C00E154B0012550C00E154B000A5F1E00E154B001CAA16034";
    defparam rom_8x4096_0_0_3.INITVAL_05 = "0x1800000000000200400001000000A8000000000E10070010021600E104B0014A90A000054B0004AA";
    defparam rom_8x4096_0_0_3.INITVAL_06 = "0x00000010080000E154B0054200000801000004A00000214000004A00000A154B0004200000000000";
    defparam rom_8x4096_0_0_3.INITVAL_07 = "0x0000001000010280000E15800004A0000EA15800004A00000E1580000A5C0000C0003001CAA160C0";
    defparam rom_8x4096_0_0_3.INITVAL_08 = "0x000000000000006040000100000000000000000801000180AC0000E05800014940000015800004AC";
    defparam rom_8x4096_0_0_3.INITVAL_09 = "0x000000000000003050090ACAA0000800455100021002A0000A174B00000000002000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_0A = "0x154A800028000000000A000000000000400000CA0000000000006000000001830000200000001000";
    defparam rom_8x4096_0_0_3.INITVAL_0B = "0x1402A000000000A10000154A800002104AA1000005400000021000A0000A0002A000080000200000";
    defparam rom_8x4096_0_0_3.INITVAL_0C = "0x12A5A000000002A0000800000100000603000000004000000000000000000000000000000A800002";
    defparam rom_8x4096_0_0_3.INITVAL_0D = "0x154AA1800212A5A0000E154AA1800E154AA1800E154AA1800212A5A0000E154AA1800E1400000002";
    defparam rom_8x4096_0_0_3.INITVAL_0E = "0x154AA180020AA560000E154AA1800E154AA1800E154AA1800E154AA180D00000000008000001000E";
    defparam rom_8x4096_0_0_3.INITVAL_0F = "0x000021800A14A55180000002A18002154AA18000000011800A1002A0000E154AA180021AA560000E";
    defparam rom_8x4096_0_0_3.INITVAL_10 = "0x00000010C00000000000000000002000000010000000014000000000000E10001100000000A1800E";
    defparam rom_8x4096_0_0_3.INITVAL_11 = "0x154AA180281140000008000800000215400000001500000000150000000A154AA180021040000000";
    defparam rom_8x4096_0_0_3.INITVAL_12 = "0x154C000002154000000E154C00000E154C000008000001000E154AA180A00000000008000800000E";
    defparam rom_8x4096_0_0_3.INITVAL_13 = "0x000800000A0AAC000000004C000002154C000000000800000A014000000C000C00000015000000EA";
    defparam rom_8x4096_0_0_3.INITVAL_14 = "0x00000000000000000000000000502000000010000000000000000000000800480000C0004C000008";
    defparam rom_8x4096_0_0_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_0_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC rom_8x4096_0_1_2 (.DIA0(scuba_vlo), .DIA1(scuba_vlo), .DIA2(scuba_vlo), 
          .DIA3(scuba_vlo), .DIA4(scuba_vlo), .DIA5(scuba_vlo), .DIA6(scuba_vlo), 
          .DIA7(scuba_vlo), .DIA8(scuba_vlo), .ADA0(scuba_vlo), .ADA1(Address_c_0), 
          .ADA2(Address_c_1), .ADA3(Address_c_2), .ADA4(Address_c_3), 
          .ADA5(Address_c_4), .ADA6(Address_c_5), .ADA7(Address_c_6), 
          .ADA8(Address_c_7), .ADA9(Address_c_8), .ADA10(Address_c_9), 
          .ADA11(Address_c_10), .ADA12(Address_c_11), .CEA(OutClockEn_c), 
          .OCEA(OutClockEn_c), .CLKA(OutClock_c), .WEA(scuba_vlo), .CSA0(scuba_vlo), 
          .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(Reset_c), .DIB0(scuba_vlo), 
          .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
          .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
          .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), .ADB3(scuba_vlo), 
          .ADB4(scuba_vlo), .ADB5(scuba_vlo), .ADB6(scuba_vlo), .ADB7(scuba_vlo), 
          .ADB8(scuba_vlo), .ADB9(scuba_vlo), .ADB10(scuba_vlo), .ADB11(scuba_vlo), 
          .ADB12(scuba_vlo), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(scuba_vlo), 
          .WEB(scuba_vlo), .CSB0(scuba_vlo), .CSB1(scuba_vlo), .CSB2(scuba_vlo), 
          .RSTB(scuba_vlo), .DOA0(Q_c_2), .DOA1(Q_c_3)) /* synthesis MEM_LPC_FILE="rom_8x4096.lpc", MEM_INIT_FILE="rom_8x4096.mem", syn_instantiated=1 */ ;
    defparam rom_8x4096_0_1_2.DATA_WIDTH_A = 2;
    defparam rom_8x4096_0_1_2.DATA_WIDTH_B = 2;
    defparam rom_8x4096_0_1_2.REGMODE_A = "NOREG";
    defparam rom_8x4096_0_1_2.REGMODE_B = "NOREG";
    defparam rom_8x4096_0_1_2.CSDECODE_A = "0b000";
    defparam rom_8x4096_0_1_2.CSDECODE_B = "0b111";
    defparam rom_8x4096_0_1_2.WRITEMODE_A = "NORMAL";
    defparam rom_8x4096_0_1_2.WRITEMODE_B = "NORMAL";
    defparam rom_8x4096_0_1_2.GSR = "ENABLED";
    defparam rom_8x4096_0_1_2.RESETMODE = "ASYNC";
    defparam rom_8x4096_0_1_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam rom_8x4096_0_1_2.INIT_DATA = "STATIC";
    defparam rom_8x4096_0_1_2.INITVAL_00 = "0x0FA4000CAA120021548000000000060BC90004DB0801D0EA74014E70A000000A4008550A00000000";
    defparam rom_8x4096_0_1_2.INITVAL_01 = "0x0600A1D4E00180C0600C0303001A550A00C000300001614000000000000C00000000000025D0A001";
    defparam rom_8x4096_0_1_2.INITVAL_02 = "0x008580600110090000C30000012280028040000400200018300600C0183000A561600C018B00180C";
    defparam rom_8x4096_0_1_2.INITVAL_03 = "0x154B001A550E00001800018200600405C300182E0600C00030018000600C01830000EB0A00C1AC30";
    defparam rom_8x4096_0_1_2.INITVAL_04 = "0x0000D0AA7001824060040583005C400600401830018000600414A2000A5A1400C00010008A60201A";
    defparam rom_8x4096_0_1_2.INITVAL_05 = "0x180000000000024074AA1580214A0006A550B80C02CB001A561400A12CA0014AD0A0051D00001800";
    defparam rom_8x4096_0_1_2.INITVAL_06 = "0x1582001A540200401800198CC0000D0BA60018CC0000C018200180C0000C01800018CC0000000004";
    defparam rom_8x4096_0_1_2.INITVAL_07 = "0x000090BA40018CC00004030001180C0004C018000180C000040180000A5C0000D0AA50008E80006A";
    defparam rom_8x4096_0_1_2.INITVAL_08 = "0x00000000000002402A590A8AA154AA054A61500D0D80002E840000A0D000014D4000071080001808";
    defparam rom_8x4096_0_1_2.INITVAL_09 = "0x054A800000000000A80C04A80180010B455000AE154EA1C0000603508000000000F00A014AA10000";
    defparam rom_8x4096_0_1_2.INITVAL_0A = "0x00001100010D00000005000000000000600000150000000002156AA00000156EA000061000212000";
    defparam rom_8x4096_0_1_2.INITVAL_0B = "0x00C401800A1540018009002811000C0028018008060580000C000801800C0C0001800E154AB10009";
    defparam rom_8x4096_0_1_2.INITVAL_0C = "0x06A581800A0001018001100090000006030000000486000068000800000A000A00000D012011000C";
    defparam rom_8x4096_0_1_2.INITVAL_0D = "0x006000800C0000018004000C01800C000C01800C000001800C000001800C000C01800401A5A1000C";
    defparam rom_8x4096_0_1_2.INITVAL_0E = "0x006001800C0000018004000A50000A154550800C0000008004004E0080C0000001800E154AA18004";
    defparam rom_8x4096_0_1_2.INITVAL_0F = "0x0B4940800002AAA1000A12A400800C000000800E154AA1800C0044018004000C01800C0600018004";
    defparam rom_8x4096_0_1_2.INITVAL_10 = "0x00000048C0000000000000000030300000001800004A50002A154AA1500C02C001800E1545008004";
    defparam rom_8x4096_0_1_2.INITVAL_11 = "0x00280000C3060C00000E154EA0000C018C00000900280000090028000009002800000C030C000000";
    defparam rom_8x4096_0_1_2.INITVAL_12 = "0x002800000C000C0000040028000004000C00000E154AA1800403000000C0000800000E154C318004";
    defparam rom_8x4096_0_1_2.INITVAL_13 = "0x15240000000B4800000A0A8400000C0000000002154E80000C060C00000D0AE4000009002800004C";
    defparam rom_8x4096_0_1_2.INITVAL_14 = "0x00000000000000000000000000061A1542A148000000000000000000000D140C00006A0A8400000D";
    defparam rom_8x4096_0_1_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_1_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC rom_8x4096_0_2_1 (.DIA0(scuba_vlo), .DIA1(scuba_vlo), .DIA2(scuba_vlo), 
          .DIA3(scuba_vlo), .DIA4(scuba_vlo), .DIA5(scuba_vlo), .DIA6(scuba_vlo), 
          .DIA7(scuba_vlo), .DIA8(scuba_vlo), .ADA0(scuba_vlo), .ADA1(Address_c_0), 
          .ADA2(Address_c_1), .ADA3(Address_c_2), .ADA4(Address_c_3), 
          .ADA5(Address_c_4), .ADA6(Address_c_5), .ADA7(Address_c_6), 
          .ADA8(Address_c_7), .ADA9(Address_c_8), .ADA10(Address_c_9), 
          .ADA11(Address_c_10), .ADA12(Address_c_11), .CEA(OutClockEn_c), 
          .OCEA(OutClockEn_c), .CLKA(OutClock_c), .WEA(scuba_vlo), .CSA0(scuba_vlo), 
          .CSA1(scuba_vlo), .CSA2(scuba_vlo), .RSTA(Reset_c), .DIB0(scuba_vlo), 
          .DIB1(scuba_vlo), .DIB2(scuba_vlo), .DIB3(scuba_vlo), .DIB4(scuba_vlo), 
          .DIB5(scuba_vlo), .DIB6(scuba_vlo), .DIB7(scuba_vlo), .DIB8(scuba_vlo), 
          .ADB0(scuba_vlo), .ADB1(scuba_vlo), .ADB2(scuba_vlo), .ADB3(scuba_vlo), 
          .ADB4(scuba_vlo), .ADB5(scuba_vlo), .ADB6(scuba_vlo), .ADB7(scuba_vlo), 
          .ADB8(scuba_vlo), .ADB9(scuba_vlo), .ADB10(scuba_vlo), .ADB11(scuba_vlo), 
          .ADB12(scuba_vlo), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(scuba_vlo), 
          .WEB(scuba_vlo), .CSB0(scuba_vlo), .CSB1(scuba_vlo), .CSB2(scuba_vlo), 
          .RSTB(scuba_vlo), .DOA0(Q_c_4), .DOA1(Q_c_5)) /* synthesis MEM_LPC_FILE="rom_8x4096.lpc", MEM_INIT_FILE="rom_8x4096.mem", syn_instantiated=1 */ ;
    defparam rom_8x4096_0_2_1.DATA_WIDTH_A = 2;
    defparam rom_8x4096_0_2_1.DATA_WIDTH_B = 2;
    defparam rom_8x4096_0_2_1.REGMODE_A = "NOREG";
    defparam rom_8x4096_0_2_1.REGMODE_B = "NOREG";
    defparam rom_8x4096_0_2_1.CSDECODE_A = "0b000";
    defparam rom_8x4096_0_2_1.CSDECODE_B = "0b111";
    defparam rom_8x4096_0_2_1.WRITEMODE_A = "NORMAL";
    defparam rom_8x4096_0_2_1.WRITEMODE_B = "NORMAL";
    defparam rom_8x4096_0_2_1.GSR = "ENABLED";
    defparam rom_8x4096_0_2_1.RESETMODE = "ASYNC";
    defparam rom_8x4096_0_2_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam rom_8x4096_0_2_1.INIT_DATA = "STATIC";
    defparam rom_8x4096_0_2_1.INITVAL_00 = "0x08200000000002400018000000000C0A80000C900A00108050000C70A00000004000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_01 = "0x020040800000251080040024000000000010AA400000000800000000000400000000000000400000";
    defparam rom_8x4096_0_2_1.INITVAL_02 = "0x00001080000320000041000090001800000000000000000255080010A24000000020010A00000250";
    defparam rom_8x4096_0_2_1.INITVAL_03 = "0x00030008000200D0AA70002700A0000005000A000A0010AA40002000A0010A24001A40000040AA40";
    defparam rom_8x4096_0_2_1.INITVAL_04 = "0x0E00000050002400A00D0824002255080000024000255080050AA7000A550A00E0000001A000E000";
    defparam rom_8x4096_0_2_1.INITVAL_05 = "0x180000000000000000000000400000020000080500010000000200400010000010A0000027000255";
    defparam rom_8x4096_0_2_1.INITVAL_06 = "0x00000000000000D0A0000C81C0000400830008500000D0AA5000814000010A00001A500000000000";
    defparam rom_8x4096_0_2_1.INITVAL_07 = "0x000040000000A0400000008001AA54000010A000002500000D0A00000A50000040000001A0C00000";
    defparam rom_8x4096_0_2_1.INITVAL_08 = "0x0000000000000180000000000000000200000804008000001C000040080000014000000380001A54";
    defparam rom_8x4096_0_2_1.INITVAL_09 = "0x080010C00000000000090D615000090AC56100061520A080050EA7A1000000001140050000000000";
    defparam rom_8x4096_0_2_1.INITVAL_0A = "0x000020800000268000000000000000006000000000000000000060000000012600000002A5400009";
    defparam rom_8x4096_0_2_1.INITVAL_0B = "0x01280180000005A180060044218006004401800E174AB10006004601800C00C801800C0000000006";
    defparam rom_8x4096_0_2_1.INITVAL_0C = "0x04A560800502C00180000309000000060300000208006000000000000005000500000600C020800C";
    defparam rom_8x4096_0_2_1.INITVAL_0D = "0x00600100061580A1800000A541800C00A5418006000020800600000180060046A0800805C5400006";
    defparam rom_8x4096_0_2_1.INITVAL_0E = "0x0060018006000020800212A001000A154FF1800C000000000E12806180150AA551800C0000018008";
    defparam rom_8x4096_0_2_1.INITVAL_0F = "0x14A681000A16A00100000ACA01000C0000010004000001800C012001800014AC0180270800208000";
    defparam rom_8x4096_0_2_1.INITVAL_10 = "0x00000000C0000000000000000018150AA550A80A1280000030000000180C0005A180040005A18008";
    defparam rom_8x4096_0_2_1.INITVAL_11 = "0x000C0000C3034C00000C000C01800C018C000006000C01000C000C000006004400000C018C000000";
    defparam rom_8x4096_0_2_1.INITVAL_12 = "0x004400000C000C000008000C00000D0AAC00000C000000000E0A2C00006A154C31800C0000000008";
    defparam rom_8x4096_0_2_1.INITVAL_13 = "0x0ACC00000A0A080000000D08000006000800000C000C00000C060C000004000C00008C000C000006";
    defparam rom_8x4096_0_2_1.INITVAL_14 = "0x00000000000000000000000000180000040000550AA550AA0A1546A1400C00CC0000010D0800000A";
    defparam rom_8x4096_0_2_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam rom_8x4096_0_2_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    OB Q_pad_7 (.I(Q_c_7), .O(Q[7]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    OB Q_pad_1 (.I(Q_c_1), .O(Q[1]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    OB Q_pad_0 (.I(Q_c_0), .O(Q[0]));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(13[23:24])
    IB Address_pad_11 (.I(Address[11]), .O(Address_c_11));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_10 (.I(Address[10]), .O(Address_c_10));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_9 (.I(Address[9]), .O(Address_c_9));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_8 (.I(Address[8]), .O(Address_c_8));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_7 (.I(Address[7]), .O(Address_c_7));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_6 (.I(Address[6]), .O(Address_c_6));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_5 (.I(Address[5]), .O(Address_c_5));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_4 (.I(Address[4]), .O(Address_c_4));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_3 (.I(Address[3]), .O(Address_c_3));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_2 (.I(Address[2]), .O(Address_c_2));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_1 (.I(Address[1]), .O(Address_c_1));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB Address_pad_0 (.I(Address[0]), .O(Address_c_0));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(9[23:30])
    IB OutClock_pad (.I(OutClock), .O(OutClock_c));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(10[16:24])
    IB OutClockEn_pad (.I(OutClockEn), .O(OutClockEn_c));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(11[16:26])
    IB Reset_pad (.I(Reset), .O(Reset_c));   // d:/codefield/verilog/diamond_design/spi_lcd/rom_8x4096.v(12[16:21])
    GSR GSR_INST (.GSR(VCC_net));
    TSALL TSALL_INST (.TSALL(scuba_vlo));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VHI i9 (.Z(VCC_net));
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

